`include "cpu_types_pkg.vh"

module branch_predictor
import cput_types_pkg::*;
(
  input logic CLK, nRST,
  input logic branck_taken,

);


